// sim/tb_fx_mul_q15.v
`timescale 1ns/1ps

module tb_fx_mul_q15;

    reg  signed [15:0] a_q15;
    reg  signed [15:0] b_q15;
    wire signed [15:0] y_q15;

    // DUT
    fx_mul_q15 dut (
        .a_q15(a_q15),
        .b_q15(b_q15),
        .y_q15(y_q15)
    );

    initial begin
        $dumpfile("tb_fx_mul_q15.vcd");
        $dumpvars(0, tb_fx_mul_q15);

        // -------------------------
        // Test 1: 0.5 * 0.5 = 0.25
        // -------------------------
        a_q15 = 16'sh4000; // 0.5
        b_q15 = 16'sh4000; // 0.5
        #10;

        // -------------------------
        // Test 2: 1.0 * 0.5 = 0.5
        // -------------------------
        a_q15 = 16'sh7FFF; // ~1.0
        b_q15 = 16'sh4000; // 0.5
        #10;

        // -------------------------
        // Test 3: -0.5 * 0.5 = -0.25
        // -------------------------
        a_q15 = -16'sh4000; // -0.5
        b_q15 =  16'sh4000; // 0.5
        #10;

        // -------------------------
        // Test 4: -0.5 * -0.5 = 0.25
        // -------------------------
        a_q15 = -16'sh4000; // -0.5
        b_q15 = -16'sh4000; // -0.5
        #10;

        // -------------------------
        // Test 5: 1.0 * 1.0 ≈ 1.0
        // -------------------------
        a_q15 = 16'sh7FFF; // ~1.0
        b_q15 = 16'sh7FFF; // ~1.0
        #10;

        #20;
        $finish;
    end

endmodule
